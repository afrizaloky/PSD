module MyXOR(a,b,x);
input a,b;
output x;

// Behavioral
assign x=a^b;

endmodule